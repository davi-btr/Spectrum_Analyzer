module VGA_interface(
	clk,
	rst_n,
	vga_clk,
	vga_blank,
	vga_sync,
	vga_R,
	vga_G,
	vga_B
);

input clk;
input rst_n;
output vga_clk;
output vga_blank;
output vga_sync;
output vga_R;
output vga_G;
output vga_B;

endmodule
