// megafunction wizard: %ALTMULT_COMPLEX%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altmult_complex 

// ============================================================
// File Name: cmplx_mult_clk.v
// Megafunction Name(s):
// 			altmult_complex
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 13.0.1 Build 232 06/12/2013 SP 1 SJ Web Edition
// ************************************************************

//Copyright (C) 1991-2013 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.

module cmplx_mult_clk (
	clock,
	dataa_imag,
	dataa_real,
	datab_imag,
	datab_real,
	result_imag,
	result_real)/* synthesis synthesis_clearbox = 1 */;

	input	  clock;
	input	[31:0]  dataa_imag;
	input	[31:0]  dataa_real;
	input	[31:0]  datab_imag;
	input	[31:0]  datab_real;
	output	[63:0]  result_imag;
	output	[63:0]  result_real;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "1"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: IMPLEMENTATION_STYLE STRING "AUTO"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
// Retrieval info: CONSTANT: PIPELINE NUMERIC "1"
// Retrieval info: CONSTANT: REPRESENTATION_A STRING "SIGNED"
// Retrieval info: CONSTANT: REPRESENTATION_B STRING "SIGNED"
// Retrieval info: CONSTANT: WIDTH_A NUMERIC "32"
// Retrieval info: CONSTANT: WIDTH_B NUMERIC "32"
// Retrieval info: CONSTANT: WIDTH_RESULT NUMERIC "64"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
// Retrieval info: USED_PORT: dataa_imag 0 0 32 0 INPUT NODEFVAL "dataa_imag[31..0]"
// Retrieval info: USED_PORT: dataa_real 0 0 32 0 INPUT NODEFVAL "dataa_real[31..0]"
// Retrieval info: USED_PORT: datab_imag 0 0 32 0 INPUT NODEFVAL "datab_imag[31..0]"
// Retrieval info: USED_PORT: datab_real 0 0 32 0 INPUT NODEFVAL "datab_real[31..0]"
// Retrieval info: USED_PORT: result_imag 0 0 64 0 OUTPUT NODEFVAL "result_imag[63..0]"
// Retrieval info: USED_PORT: result_real 0 0 64 0 OUTPUT NODEFVAL "result_real[63..0]"
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: @dataa_imag 0 0 32 0 dataa_imag 0 0 32 0
// Retrieval info: CONNECT: @dataa_real 0 0 32 0 dataa_real 0 0 32 0
// Retrieval info: CONNECT: @datab_imag 0 0 32 0 datab_imag 0 0 32 0
// Retrieval info: CONNECT: @datab_real 0 0 32 0 datab_real 0 0 32 0
// Retrieval info: CONNECT: result_imag 0 0 64 0 @result_imag 0 0 64 0
// Retrieval info: CONNECT: result_real 0 0 64 0 @result_real 0 0 64 0
// Retrieval info: GEN_FILE: TYPE_NORMAL cmplx_mult_clk.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL cmplx_mult_clk.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL cmplx_mult_clk.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL cmplx_mult_clk.bsf TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL cmplx_mult_clk_inst.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL cmplx_mult_clk_bb.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL cmplx_mult_clk_syn.v TRUE
// Retrieval info: LIB_FILE: altera_mf
